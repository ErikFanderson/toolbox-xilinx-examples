//==============================================================================
// Author: Erik Anderson 
// Email: efa@eecs.berkeley.edu 
// Description: <Insert Description Here> 
// Naming conventions:
//    signals => snake_case
//    Parameters (aliasing signal values) => SNAKE_CASE with all caps
//    Parameters (not aliasing signal values) => CamelCase 
//==============================================================================
`timescale 1ns/1ps
`default_nettype none

interface led_blink_bfm;
//-----------------------------------------------------------------------------
// Imports and macros 
//-----------------------------------------------------------------------------
import uvm_pkg::*;
import led_blink_pkg::*;
`include "uvm_macros.svh"
//-----------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Parameters 
//------------------------------------------------------------------------------
// Interface/Simulation Parameters
parameter real ClockCycle = 1.0;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Constants (localparam) 
//------------------------------------------------------------------------------
// Interface/Simulation constants 
localparam real HalfClockCycle = ClockCycle/2.0;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Inputs/Outputs 
//------------------------------------------------------------------------------
logic clk_p;
logic clk_n;
logic led;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Initial stuff
//------------------------------------------------------------------------------
initial begin
    clk_p = 0;
    clk_n = 1;
    forever begin
        #(HalfClockCycle);
        clk_p = ~clk_p;
        clk_n = ~clk_n;
    end
end
//------------------------------------------------------------------------------
endinterface : led_blink_bfm 

`default_nettype wire 
