//==============================================================================
// Author: Erik Anderson 
// Email: efa@eecs.berkeley.edu 
// Description: <Insert Description Here> 
// Naming conventions:
//    signals => snake_case
//    Parameters (aliasing signal values) => SNAKE_CASE with all caps
//    Parameters (not aliasing signal values) => CamelCase 
//==============================================================================
`timescale 1ns/1ps
`default_nettype none

interface led_blink_bfm;
//-----------------------------------------------------------------------------
// Imports and macros 
//-----------------------------------------------------------------------------
import uvm_pkg::*;
import led_blink_pkg::*;
`include "uvm_macros.svh"
//-----------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Parameters 
//------------------------------------------------------------------------------
// Interface/Simulation Parameters
parameter real ClockCycle = 1.0;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Constants (localparam) 
//------------------------------------------------------------------------------
// Interface/Simulation constants 
localparam real HalfClockCycle = ClockCycle/2.0;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Inputs/Outputs 
//------------------------------------------------------------------------------
logic i_clk;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Initial stuff
//------------------------------------------------------------------------------
initial begin
    i_clk = 0;
    forever begin
        #(HalfClockCycle);
        i_clk = ~i_clk;
    end
end
//------------------------------------------------------------------------------
endinterface : led_blink_bfm 

`default_nettype wire 
